parameter N = 3;