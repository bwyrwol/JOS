module test(input a, output y);

assign y = a;

endmodule
